library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.std_logic_misc.ALL;
use ieee.math_real.all;
Library IEEE_PROPOSED;
Use IEEE_PROPOSED.FIXED_PKG.All;

package ZCONSTANTS is    

    constant ZN12 : integer := -12;
    constant ZN11 : integer := -11;
    constant ZN10 : integer := -10;
    constant ZN9 : integer := -9;
    constant ZN8 : integer := -8;
    constant ZN7 : integer := -7;
    constant ZN6 : integer := -6;
    constant ZN5 : integer := -5;
    constant ZN4 : integer := -4;
    constant ZN3 : integer := -3;
    constant ZN2 : integer := -2;
    constant ZN1 : integer := -1;
    constant Z00 : integer := 0;
    constant Z01 : integer := 1;
    constant Z02 : integer := 2;
    constant Z03 : integer := 3;
    constant Z04 : integer := 4;
    constant Z05 : integer := 5;    
    constant Z06 : integer := 6;
    constant Z07 : integer := 7;
    constant Z08 : integer := 8;
    constant Z09 : integer := 9;
    constant Z10 : integer := 10;
    constant Z11 : integer := 11;
    constant Z12 : integer := 12;
    constant Z13 : integer := 13;
    constant Z14 : integer := 14;
    constant Z15 : integer := 15;    
    constant Z16 : integer := 16;
    constant Z17 : integer := 17;
    constant Z18 : integer := 18;
    constant Z19 : integer := 19;
    constant Z20 : integer := 20;
    constant Z21 : integer := 21;
    constant Z22 : integer := 22;
    constant Z23 : integer := 23;   
    constant Z24 : integer := 24;      
    constant Z25 : integer := 25;    
    constant Z26 : integer := 26;
    constant Z27 : integer := 27;
    constant Z28 : integer := 28;
    constant Z29 : integer := 29;     
    constant Z30 : integer := 30;
    constant Z31 : integer := 31;
    constant Z32 : integer := 32;
    constant Z33 : integer := 33;
    constant Z34 : integer := 34;
    constant Z35 : integer := 35;    
    constant Z36 : integer := 36;
    constant Z37 : integer := 37;
    constant Z38 : integer := 38;
    constant Z39 : integer := 39;
    constant Z40 : integer := 40;
    constant Z41 : integer := 41;
    constant Z42 : integer := 42;
    constant Z43 : integer := 43;
    constant Z44 : integer := 44;
    constant Z45 : integer := 45;    
    constant Z46 : integer := 46;
    constant Z47 : integer := 47;
    constant Z48 : integer := 48;
    constant Z49 : integer := 49;
    constant Z50 : integer := 50;   
    constant Z51 : integer := 51;
    constant Z52 : integer := 52;
    constant Z53 : integer := 53;
    constant Z54 : integer := 54;
    constant Z55 : integer := 55;    
    constant Z56 : integer := 56;
    constant Z57 : integer := 57;
    constant Z58 : integer := 58;
    constant Z59 : integer := 59;
    constant Z60 : integer := 60;   
    constant Z61 : integer := 61;
    constant Z62 : integer := 62;
    constant Z63 : integer := 63;
    constant Z64 : integer := 64;
    constant Z65 : integer := 65;
    constant Z66 : integer := 66;
    constant Z67 : integer := 67;
    constant Z68 : integer := 68;
    constant Z69 : integer := 69;
            
    constant YN12 : integer := -12;
    constant YN11 : integer := -11;
    constant YN10 : integer := -10;
    constant YN9 : integer := -9;
    constant YN8 : integer := -8;
    constant YN7 : integer := -7;
    constant YN6 : integer := -6;
    constant YN5 : integer := -5;
    constant YN4 : integer := -4;
    constant YN3 : integer := -3;
    constant YN2 : integer := -2;
    constant YN1 : integer := -1;
    constant Y00 : integer := 0;
    constant Y01 : integer := 1;
    constant Y02 : integer := 2;
    constant Y03 : integer := 3;
    constant Y04 : integer := 4;
    constant Y05 : integer := 5;    
    constant Y06 : integer := 6;
    constant Y07 : integer := 7;
    constant Y08 : integer := 8;
    constant Y09 : integer := 9;
    constant Y10 : integer := 10;
    constant Y11 : integer := 11;
    constant Y12 : integer := 12;
    constant Y13 : integer := 13;
    constant Y14 : integer := 14;
    constant Y15 : integer := 15;    
    constant Y16 : integer := 16;
    constant Y17 : integer := 17;
    constant Y18 : integer := 18;
    constant Y19 : integer := 19;
    constant Y20 : integer := 20;
    constant Y21 : integer := 21;
    constant Y22 : integer := 22;
    constant Y23 : integer := 23;   
    constant Y24 : integer := 24;      
    constant Y25 : integer := 25;    
    constant Y26 : integer := 26;
    constant Y27 : integer := 27;
    constant Y28 : integer := 28;
    constant Y29 : integer := 29;     
    constant Y30 : integer := 30;
    constant Y31 : integer := 31;
    constant Y32 : integer := 32;
    constant Y33 : integer := 33;
    constant Y34 : integer := 34;
    constant Y35 : integer := 35;    
    constant Y36 : integer := 36;
    constant Y37 : integer := 37;
    constant Y38 : integer := 38;
    constant Y39 : integer := 39;
    constant Y40 : integer := 40;
    constant Y41 : integer := 41;
    constant Y42 : integer := 42;
    constant Y43 : integer := 43;
    constant Y44 : integer := 44;
    constant Y45 : integer := 45;    
    constant Y46 : integer := 46;
    constant Y47 : integer := 47;
    constant Y48 : integer := 48;
    constant Y49 : integer := 49;
    constant Y50 : integer := 50;   
    constant Y51 : integer := 51;
    constant Y52 : integer := 52;
    constant Y53 : integer := 53;
    constant Y54 : integer := 54;
    constant Y55 : integer := 55;    
    constant Y56 : integer := 56;
    constant Y57 : integer := 57;
    constant Y58 : integer := 58;
    constant Y59 : integer := 59;
    constant Y60 : integer := 60;   
    constant Y61 : integer := 61;
    constant Y62 : integer := 62;
    constant Y63 : integer := 63;
    constant Y64 : integer := 64;
    constant Y65 : integer := 65;
    constant Y66 : integer := 66;
    constant Y67 : integer := 67;
    constant Y68 : integer := 68;
    constant Y69 : integer := 69;
    
    constant SN12 : integer := -12;
    constant SN11 : integer := -11;
    constant SN10 : integer := -10;
    constant SN9 : integer := -9;
    constant SN8 : integer := -8;
    constant SN7 : integer := -7;
    constant SN6 : integer := -6;
    constant SN5 : integer := -5;
    constant SN4 : integer := -4;
    constant SN3 : integer := -3;
    constant SN2 : integer := -2;
    constant SN1 : integer := -1;
    constant S00 : integer := 0;
    constant S01 : integer := 1;
    constant S02 : integer := 2;
    constant S03 : integer := 3;
    constant S04 : integer := 4;
    constant S05 : integer := 5;    
    constant S06 : integer := 6;
    constant S07 : integer := 7;
    constant S08 : integer := 8;
    constant S09 : integer := 9;
    constant S10 : integer := 10;
    constant S11 : integer := 11;
    constant S12 : integer := 12;
    constant S13 : integer := 13;
    constant S14 : integer := 14;
    constant S15 : integer := 15;    
    constant S16 : integer := 16;
    constant S17 : integer := 17;
    constant S18 : integer := 18;
    constant S19 : integer := 19;
    constant S20 : integer := 20;
    constant S21 : integer := 21;
    constant S22 : integer := 22;
    constant S23 : integer := 23;   
    constant S24 : integer := 24;      
    constant S25 : integer := 25;    
    constant S26 : integer := 26;
    constant S27 : integer := 27;
    constant S28 : integer := 28;
    constant S29 : integer := 29;     
    constant S30 : integer := 30;
    constant S31 : integer := 31;
    constant S32 : integer := 32;
    constant S33 : integer := 33;
    constant S34 : integer := 34;
    constant S35 : integer := 35;    
    constant S36 : integer := 36;
    constant S37 : integer := 37;
    constant S38 : integer := 38;
    constant S39 : integer := 39;
    constant S40 : integer := 40;
    constant S41 : integer := 41;
    constant S42 : integer := 42;
    constant S43 : integer := 43;
    constant S44 : integer := 44;
    constant S45 : integer := 45;    
    constant S46 : integer := 46;
    constant S47 : integer := 47;
    constant S48 : integer := 48;
    constant S49 : integer := 49;
    constant S50 : integer := 50;   
    constant S51 : integer := 51;
    constant S52 : integer := 52;
    constant S53 : integer := 53;
    constant S54 : integer := 54;
    constant S55 : integer := 55;    
    constant S56 : integer := 56;
    constant S57 : integer := 57;
    constant S58 : integer := 58;
    constant S59 : integer := 59;
    constant S60 : integer := 60;   
    constant S61 : integer := 61;
    constant S62 : integer := 62;
    constant S63 : integer := 63;
    constant S64 : integer := 64;
    constant S65 : integer := 65;
    constant S66 : integer := 66;
    constant S67 : integer := 67;
    constant S68 : integer := 68;
    constant S69 : integer := 69;
    
end ZCONSTANTS;
